`timescale 1ps/1ps

module p5_tb;
    reg [2:0] a;
    reg [2:0] b;
    wire [5:0] f;

    p5 mult(a,b,f);

    always
    begin
        $dumpfile("p5.vcd");
        $dumpvars(0,p5_tb);

        a = 0;
        b = 0;
        #10
        b = 1;
        #10
        b = 2;
        #10
        b = 3;
        #10
        b = 4;
        #10
        b = 5;
        #10
        b = 6;
        #10
        b = 7;
        #10

        a = 1;
        b = 0;
        #10
        b = 1;
        #10
        b = 2;
        #10
        b = 3;
        #10
        b = 4;
        #10
        b = 5;
        #10
        b = 6;
        #10
        b = 7;
        #10

        a = 2;
        b = 0;
        #10
        b = 1;
        #10
        b = 2;
        #10
        b = 3;
        #10
        b = 4;
        #10
        b = 5;
        #10
        b = 6;
        #10
        b = 7;
        #10

        a = 3;
        b = 0;
        #10
        b = 1;
        #10
        b = 2;
        #10
        b = 3;
        #10
        b = 4;
        #10
        b = 5;
        #10
        b = 6;
        #10
        b = 7;
        #10

        a = 4;
        b = 0;
        #10
        b = 1;
        #10
        b = 2;
        #10
        b = 3;
        #10
        b = 4;
        #10
        b = 5;
        #10
        b = 6;
        #10
        b = 7;
        #10

        a = 5;
        b = 0;
        #10
        b = 1;
        #10
        b = 2;
        #10
        b = 3;
        #10
        b = 4;
        #10
        b = 5;
        #10
        b = 6;
        #10
        b = 7;
        #10

        a = 6;
        b = 0;
        #10
        b = 1;
        #10
        b = 2;
        #10
        b = 3;
        #10
        b = 4;
        #10
        b = 5;
        #10
        b = 6;
        #10
        b = 7;
        #10

        a = 7;
        b = 0;
        #10
        b = 1;
        #10
        b = 2;
        #10
        b = 3;
        #10
        b = 4;
        #10
        b = 5;
        #10
        b = 6;
        #10
        b = 7;
        #10

        $finish;
    end
endmodule